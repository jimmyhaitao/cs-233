module blackbox(l, s, i, w);
    output l;
    input  s, i, w;
    wire   w01, w07, w08, w15, w25, w31, w33, w42, w48, w49, w52, w58, w60, w63, w64, w67, w72, w80, w82, w85, w91, w92, w96;
    or  o88(l, w63, w92, w80);
    and a79(w63, w52, w60, w48);
    not n93(w48, w25);
    and a78(w92, w60, w25, w52);
    and a90(w80, w01, w07);
    not n53(w01, w60);
    or  o26(w07, w15, w58);
    and a43(w15, w52, w25);
    and a68(w58, w42, w52);
    not n81(w42, w25);
    and a65(w60, i, w82);
    or  o94(w82, w, s);
    and a71(w25, w67, w31);
    not n4(w67, s);
    or  o35(w31, w85, w72);
    not n21(w85, w);
    and a3(w72, i, w33);
    not n62(w33, i);
    or  o41(w52, w08, w96);
    and a97(w08, w64, w49);
    not n61(w64, i);
    not n5(w49, s);
    and a34(w96, w91, w, i);
    not n18(w91, s);
endmodule // blackbox
